class transaction;
rand bit d;
  bit q;
endclass
