interface intf(input logic clk,reset);
  logic d;
  logic q;
endinterface
