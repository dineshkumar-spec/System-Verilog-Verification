interface intf;
  logic a,b,c;
  logic sum,cout;
endinterface
